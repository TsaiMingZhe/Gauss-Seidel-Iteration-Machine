module testbench (
    ports
);
    
endmodule